-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb5",
     9 => x"d4080b0b",
    10 => x"0bb5d808",
    11 => x"0b0b0bb5",
    12 => x"dc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b5dc0c0b",
    16 => x"0b0bb5d8",
    17 => x"0c0b0b0b",
    18 => x"b5d40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0baf84",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b5d47080",
    57 => x"c084278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188fe04",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb5e40c",
    65 => x"9f0bb5e8",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b5e808ff",
    69 => x"05b5e80c",
    70 => x"b5e80880",
    71 => x"25eb38b5",
    72 => x"e408ff05",
    73 => x"b5e40cb5",
    74 => x"e4088025",
    75 => x"d738800b",
    76 => x"b5e80c80",
    77 => x"0bb5e40c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb5e408",
    97 => x"258f3882",
    98 => x"bd2db5e4",
    99 => x"08ff05b5",
   100 => x"e40c82ff",
   101 => x"04b5e408",
   102 => x"b5e80853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b5e408a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b5e8",
   111 => x"088105b5",
   112 => x"e80cb5e8",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb5e80c",
   116 => x"b5e40881",
   117 => x"05b5e40c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b5",
   122 => x"e8088105",
   123 => x"b5e80cb5",
   124 => x"e808a02e",
   125 => x"0981068e",
   126 => x"38800bb5",
   127 => x"e80cb5e4",
   128 => x"088105b5",
   129 => x"e40c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb5ec",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb5ec0c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b5",
   169 => x"ec088407",
   170 => x"b5ec0c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb29c",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b5ec0852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b5d40c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c8da32d",
   216 => x"0284050d",
   217 => x"0402fc05",
   218 => x"0dec5192",
   219 => x"710c86a4",
   220 => x"2d82710c",
   221 => x"0284050d",
   222 => x"0402fc05",
   223 => x"0d8da32d",
   224 => x"ec5180c2",
   225 => x"710c86a4",
   226 => x"2d80710c",
   227 => x"0284050d",
   228 => x"0402d005",
   229 => x"0d7d5480",
   230 => x"5ba40bec",
   231 => x"0c7352b5",
   232 => x"f051a6c2",
   233 => x"2db5d408",
   234 => x"7b2e81ab",
   235 => x"38b5f408",
   236 => x"70f80c89",
   237 => x"1580f52d",
   238 => x"8a1680f5",
   239 => x"2d718280",
   240 => x"29058817",
   241 => x"80f52d70",
   242 => x"84808029",
   243 => x"12f40c7e",
   244 => x"ff155c5e",
   245 => x"57555658",
   246 => x"767b2e8b",
   247 => x"38811a77",
   248 => x"812a585a",
   249 => x"76f738f7",
   250 => x"1a5a815b",
   251 => x"80782580",
   252 => x"e6387952",
   253 => x"7651848b",
   254 => x"2db6bc52",
   255 => x"b5f051a8",
   256 => x"f82db5d4",
   257 => x"08802eb8",
   258 => x"38b6bc5c",
   259 => x"83fc597b",
   260 => x"7084055d",
   261 => x"087081ff",
   262 => x"0671882a",
   263 => x"7081ff06",
   264 => x"73902a70",
   265 => x"81ff0675",
   266 => x"982ae80c",
   267 => x"e80c58e8",
   268 => x"0c57e80c",
   269 => x"fc1a5a53",
   270 => x"788025d3",
   271 => x"3888c704",
   272 => x"b5d4085b",
   273 => x"848058b5",
   274 => x"f051a8cb",
   275 => x"2dfc8018",
   276 => x"81185858",
   277 => x"87ec0486",
   278 => x"b72d800b",
   279 => x"ec0c7a80",
   280 => x"2e8d38b2",
   281 => x"a0518fa0",
   282 => x"2d8da32d",
   283 => x"88f504b3",
   284 => x"a4518fa0",
   285 => x"2d7ab5d4",
   286 => x"0c02b005",
   287 => x"0d0402f4",
   288 => x"050d850b",
   289 => x"ec0c8d84",
   290 => x"2d89ee2d",
   291 => x"81f82d9d",
   292 => x"df2db5d4",
   293 => x"08802e80",
   294 => x"c0388791",
   295 => x"51aeff2d",
   296 => x"b2a0518f",
   297 => x"a02d8da3",
   298 => x"2d89fa2d",
   299 => x"8fb02db2",
   300 => x"e40b80f5",
   301 => x"2d70822b",
   302 => x"8406b2d8",
   303 => x"0b80f52d",
   304 => x"83067107",
   305 => x"fc0c5353",
   306 => x"8652b5d4",
   307 => x"088538b5",
   308 => x"d4085271",
   309 => x"ec0c89a9",
   310 => x"04800bb5",
   311 => x"d40c028c",
   312 => x"050d0471",
   313 => x"980c04ff",
   314 => x"b008b5d4",
   315 => x"0c04810b",
   316 => x"ffb00c04",
   317 => x"800bffb0",
   318 => x"0c0402f4",
   319 => x"050d8afc",
   320 => x"04b5d408",
   321 => x"81f02e09",
   322 => x"81068938",
   323 => x"810bb488",
   324 => x"0c8afc04",
   325 => x"b5d40881",
   326 => x"e02e0981",
   327 => x"06893881",
   328 => x"0bb48c0c",
   329 => x"8afc04b5",
   330 => x"d40852b4",
   331 => x"8c08802e",
   332 => x"8838b5d4",
   333 => x"08818005",
   334 => x"5271842c",
   335 => x"728f0653",
   336 => x"53b48808",
   337 => x"802e9938",
   338 => x"728429b3",
   339 => x"c8057213",
   340 => x"81712b70",
   341 => x"09730806",
   342 => x"730c5153",
   343 => x"538af204",
   344 => x"728429b3",
   345 => x"c8057213",
   346 => x"83712b72",
   347 => x"0807720c",
   348 => x"5353800b",
   349 => x"b48c0c80",
   350 => x"0bb4880c",
   351 => x"b5fc518b",
   352 => x"fd2db5d4",
   353 => x"08ff24fe",
   354 => x"f838800b",
   355 => x"b5d40c02",
   356 => x"8c050d04",
   357 => x"02f8050d",
   358 => x"b3c8528f",
   359 => x"51807270",
   360 => x"8405540c",
   361 => x"ff115170",
   362 => x"8025f238",
   363 => x"0288050d",
   364 => x"0402f005",
   365 => x"0d755189",
   366 => x"f42d7082",
   367 => x"2cfc06b3",
   368 => x"c8117210",
   369 => x"9e067108",
   370 => x"70722a70",
   371 => x"83068274",
   372 => x"2b700974",
   373 => x"06760c54",
   374 => x"51565753",
   375 => x"515389ee",
   376 => x"2d71b5d4",
   377 => x"0c029005",
   378 => x"0d0402fc",
   379 => x"050d7251",
   380 => x"80710c80",
   381 => x"0b84120c",
   382 => x"0284050d",
   383 => x"0402f005",
   384 => x"0d757008",
   385 => x"84120853",
   386 => x"5353ff54",
   387 => x"71712ea8",
   388 => x"3889f42d",
   389 => x"84130870",
   390 => x"84291488",
   391 => x"11700870",
   392 => x"81ff0684",
   393 => x"18088111",
   394 => x"8706841a",
   395 => x"0c535155",
   396 => x"51515189",
   397 => x"ee2d7154",
   398 => x"73b5d40c",
   399 => x"0290050d",
   400 => x"0402f805",
   401 => x"0d89f42d",
   402 => x"e008708b",
   403 => x"2a708106",
   404 => x"51525270",
   405 => x"802e9d38",
   406 => x"b5fc0870",
   407 => x"8429b684",
   408 => x"057381ff",
   409 => x"06710c51",
   410 => x"51b5fc08",
   411 => x"81118706",
   412 => x"b5fc0c51",
   413 => x"800bb6a4",
   414 => x"0c89e72d",
   415 => x"89ee2d02",
   416 => x"88050d04",
   417 => x"02fc050d",
   418 => x"b5fc518b",
   419 => x"ea2d8b94",
   420 => x"2d8cc151",
   421 => x"89e32d02",
   422 => x"84050d04",
   423 => x"b6a808b5",
   424 => x"d40c0402",
   425 => x"fc050d8d",
   426 => x"ad0489fa",
   427 => x"2d80f651",
   428 => x"8bb12db5",
   429 => x"d408f338",
   430 => x"80da518b",
   431 => x"b12db5d4",
   432 => x"08e838b5",
   433 => x"d408b494",
   434 => x"0cb5d408",
   435 => x"5184f02d",
   436 => x"0284050d",
   437 => x"0402ec05",
   438 => x"0d765480",
   439 => x"52870b88",
   440 => x"1580f52d",
   441 => x"56537472",
   442 => x"248338a0",
   443 => x"53725182",
   444 => x"f92d8112",
   445 => x"8b1580f5",
   446 => x"2d545272",
   447 => x"7225de38",
   448 => x"0294050d",
   449 => x"0402f005",
   450 => x"0db6a808",
   451 => x"5481f82d",
   452 => x"800bb6ac",
   453 => x"0c730880",
   454 => x"2e818038",
   455 => x"820bb5e8",
   456 => x"0cb6ac08",
   457 => x"8f06b5e4",
   458 => x"0c730852",
   459 => x"71832e96",
   460 => x"38718326",
   461 => x"89387181",
   462 => x"2eaf388f",
   463 => x"86047185",
   464 => x"2e9f388f",
   465 => x"86048814",
   466 => x"80f52d84",
   467 => x"1508b0e8",
   468 => x"53545285",
   469 => x"fe2d7184",
   470 => x"29137008",
   471 => x"52528f8a",
   472 => x"0473518d",
   473 => x"d52d8f86",
   474 => x"04b49008",
   475 => x"8815082c",
   476 => x"70810651",
   477 => x"5271802e",
   478 => x"8738b0ec",
   479 => x"518f8304",
   480 => x"b0f05185",
   481 => x"fe2d8414",
   482 => x"085185fe",
   483 => x"2db6ac08",
   484 => x"8105b6ac",
   485 => x"0c8c1454",
   486 => x"8e950402",
   487 => x"90050d04",
   488 => x"71b6a80c",
   489 => x"8e852db6",
   490 => x"ac08ff05",
   491 => x"b6b00c04",
   492 => x"02e8050d",
   493 => x"b6a808b6",
   494 => x"b4085755",
   495 => x"87518bb1",
   496 => x"2db5d408",
   497 => x"812a7081",
   498 => x"06515271",
   499 => x"802ea038",
   500 => x"8fd60489",
   501 => x"fa2d8751",
   502 => x"8bb12db5",
   503 => x"d408f438",
   504 => x"b4940881",
   505 => x"3270b494",
   506 => x"0c705252",
   507 => x"84f02d80",
   508 => x"fe518bb1",
   509 => x"2db5d408",
   510 => x"802ea638",
   511 => x"b4940880",
   512 => x"2e913880",
   513 => x"0bb4940c",
   514 => x"805184f0",
   515 => x"2d909304",
   516 => x"89fa2d80",
   517 => x"fe518bb1",
   518 => x"2db5d408",
   519 => x"f33886e5",
   520 => x"2db49408",
   521 => x"903881fd",
   522 => x"518bb12d",
   523 => x"81fa518b",
   524 => x"b12d95e6",
   525 => x"0481f551",
   526 => x"8bb12db5",
   527 => x"d408812a",
   528 => x"70810651",
   529 => x"5271802e",
   530 => x"af38b6b0",
   531 => x"08527180",
   532 => x"2e8938ff",
   533 => x"12b6b00c",
   534 => x"90f804b6",
   535 => x"ac0810b6",
   536 => x"ac080570",
   537 => x"84291651",
   538 => x"52881208",
   539 => x"802e8938",
   540 => x"ff518812",
   541 => x"0852712d",
   542 => x"81f2518b",
   543 => x"b12db5d4",
   544 => x"08812a70",
   545 => x"81065152",
   546 => x"71802eb1",
   547 => x"38b6ac08",
   548 => x"ff11b6b0",
   549 => x"08565353",
   550 => x"73722589",
   551 => x"388114b6",
   552 => x"b00c91bd",
   553 => x"04721013",
   554 => x"70842916",
   555 => x"51528812",
   556 => x"08802e89",
   557 => x"38fe5188",
   558 => x"12085271",
   559 => x"2d81fd51",
   560 => x"8bb12db5",
   561 => x"d408812a",
   562 => x"70810651",
   563 => x"5271802e",
   564 => x"ad38b6b0",
   565 => x"08802e89",
   566 => x"38800bb6",
   567 => x"b00c91fe",
   568 => x"04b6ac08",
   569 => x"10b6ac08",
   570 => x"05708429",
   571 => x"16515288",
   572 => x"1208802e",
   573 => x"8938fd51",
   574 => x"88120852",
   575 => x"712d81fa",
   576 => x"518bb12d",
   577 => x"b5d40881",
   578 => x"2a708106",
   579 => x"51527180",
   580 => x"2eae38b6",
   581 => x"ac08ff11",
   582 => x"5452b6b0",
   583 => x"08732588",
   584 => x"3872b6b0",
   585 => x"0c92c004",
   586 => x"71101270",
   587 => x"84291651",
   588 => x"52881208",
   589 => x"802e8938",
   590 => x"fc518812",
   591 => x"0852712d",
   592 => x"b6b00870",
   593 => x"53547380",
   594 => x"2e8a388c",
   595 => x"15ff1555",
   596 => x"5592c604",
   597 => x"820bb5e8",
   598 => x"0c718f06",
   599 => x"b5e40c81",
   600 => x"eb518bb1",
   601 => x"2db5d408",
   602 => x"812a7081",
   603 => x"06515271",
   604 => x"802ead38",
   605 => x"7408852e",
   606 => x"098106a4",
   607 => x"38881580",
   608 => x"f52dff05",
   609 => x"52718816",
   610 => x"81b72d71",
   611 => x"982b5271",
   612 => x"80258838",
   613 => x"800b8816",
   614 => x"81b72d74",
   615 => x"518dd52d",
   616 => x"81f4518b",
   617 => x"b12db5d4",
   618 => x"08812a70",
   619 => x"81065152",
   620 => x"71802eb3",
   621 => x"38740885",
   622 => x"2e098106",
   623 => x"aa388815",
   624 => x"80f52d81",
   625 => x"05527188",
   626 => x"1681b72d",
   627 => x"7181ff06",
   628 => x"8b1680f5",
   629 => x"2d545272",
   630 => x"72278738",
   631 => x"72881681",
   632 => x"b72d7451",
   633 => x"8dd52d80",
   634 => x"da518bb1",
   635 => x"2db5d408",
   636 => x"812a7081",
   637 => x"06515271",
   638 => x"802e81a6",
   639 => x"38b6a808",
   640 => x"b6b00855",
   641 => x"5373802e",
   642 => x"8a388c13",
   643 => x"ff155553",
   644 => x"94850472",
   645 => x"08527182",
   646 => x"2ea63871",
   647 => x"82268938",
   648 => x"71812ea9",
   649 => x"3895a204",
   650 => x"71832eb1",
   651 => x"3871842e",
   652 => x"09810680",
   653 => x"ed388813",
   654 => x"08518fa0",
   655 => x"2d95a204",
   656 => x"b6b00851",
   657 => x"88130852",
   658 => x"712d95a2",
   659 => x"04810b88",
   660 => x"14082bb4",
   661 => x"900832b4",
   662 => x"900c94f8",
   663 => x"04881380",
   664 => x"f52d8105",
   665 => x"8b1480f5",
   666 => x"2d535471",
   667 => x"74248338",
   668 => x"80547388",
   669 => x"1481b72d",
   670 => x"8e852d95",
   671 => x"a2047508",
   672 => x"802ea238",
   673 => x"7508518b",
   674 => x"b12db5d4",
   675 => x"08810652",
   676 => x"71802e8b",
   677 => x"38b6b008",
   678 => x"51841608",
   679 => x"52712d88",
   680 => x"165675da",
   681 => x"38805480",
   682 => x"0bb5e80c",
   683 => x"738f06b5",
   684 => x"e40ca052",
   685 => x"73b6b008",
   686 => x"2e098106",
   687 => x"9838b6ac",
   688 => x"08ff0574",
   689 => x"32700981",
   690 => x"05707207",
   691 => x"9f2a9171",
   692 => x"31515153",
   693 => x"53715182",
   694 => x"f92d8114",
   695 => x"548e7425",
   696 => x"c638b494",
   697 => x"085271b5",
   698 => x"d40c0298",
   699 => x"050d0402",
   700 => x"f4050dd4",
   701 => x"5281ff72",
   702 => x"0c710853",
   703 => x"81ff720c",
   704 => x"72882b83",
   705 => x"fe800672",
   706 => x"087081ff",
   707 => x"06515253",
   708 => x"81ff720c",
   709 => x"72710788",
   710 => x"2b720870",
   711 => x"81ff0651",
   712 => x"525381ff",
   713 => x"720c7271",
   714 => x"07882b72",
   715 => x"087081ff",
   716 => x"067207b5",
   717 => x"d40c5253",
   718 => x"028c050d",
   719 => x"0402f405",
   720 => x"0d747671",
   721 => x"81ff06d4",
   722 => x"0c5353b6",
   723 => x"b8088538",
   724 => x"71892b52",
   725 => x"71982ad4",
   726 => x"0c71902a",
   727 => x"7081ff06",
   728 => x"d40c5171",
   729 => x"882a7081",
   730 => x"ff06d40c",
   731 => x"517181ff",
   732 => x"06d40c72",
   733 => x"902a7081",
   734 => x"ff06d40c",
   735 => x"51d40870",
   736 => x"81ff0651",
   737 => x"5182b8bf",
   738 => x"527081ff",
   739 => x"2e098106",
   740 => x"943881ff",
   741 => x"0bd40cd4",
   742 => x"087081ff",
   743 => x"06ff1454",
   744 => x"515171e5",
   745 => x"3870b5d4",
   746 => x"0c028c05",
   747 => x"0d0402fc",
   748 => x"050d81c7",
   749 => x"5181ff0b",
   750 => x"d40cff11",
   751 => x"51708025",
   752 => x"f4380284",
   753 => x"050d0402",
   754 => x"f4050d81",
   755 => x"ff0bd40c",
   756 => x"93538052",
   757 => x"87fc80c1",
   758 => x"5196bd2d",
   759 => x"b5d4088b",
   760 => x"3881ff0b",
   761 => x"d40c8153",
   762 => x"97f40497",
   763 => x"ae2dff13",
   764 => x"5372df38",
   765 => x"72b5d40c",
   766 => x"028c050d",
   767 => x"0402ec05",
   768 => x"0d810bb6",
   769 => x"b80c8454",
   770 => x"d008708f",
   771 => x"2a708106",
   772 => x"51515372",
   773 => x"f33872d0",
   774 => x"0c97ae2d",
   775 => x"b0f45185",
   776 => x"fe2dd008",
   777 => x"708f2a70",
   778 => x"81065151",
   779 => x"5372f338",
   780 => x"810bd00c",
   781 => x"b1538052",
   782 => x"84d480c0",
   783 => x"5196bd2d",
   784 => x"b5d40881",
   785 => x"2e933872",
   786 => x"822ebd38",
   787 => x"ff135372",
   788 => x"e538ff14",
   789 => x"5473ffb0",
   790 => x"3897ae2d",
   791 => x"83aa5284",
   792 => x"9c80c851",
   793 => x"96bd2db5",
   794 => x"d408812e",
   795 => x"09810692",
   796 => x"3895ef2d",
   797 => x"b5d40883",
   798 => x"ffff0653",
   799 => x"7283aa2e",
   800 => x"9d3897c7",
   801 => x"2d999904",
   802 => x"b1805185",
   803 => x"fe2d8053",
   804 => x"9ae704b1",
   805 => x"985185fe",
   806 => x"2d80549a",
   807 => x"b90481ff",
   808 => x"0bd40cb1",
   809 => x"5497ae2d",
   810 => x"8fcf5380",
   811 => x"5287fc80",
   812 => x"f75196bd",
   813 => x"2db5d408",
   814 => x"55b5d408",
   815 => x"812e0981",
   816 => x"069b3881",
   817 => x"ff0bd40c",
   818 => x"820a5284",
   819 => x"9c80e951",
   820 => x"96bd2db5",
   821 => x"d408802e",
   822 => x"8d3897ae",
   823 => x"2dff1353",
   824 => x"72c9389a",
   825 => x"ac0481ff",
   826 => x"0bd40cb5",
   827 => x"d4085287",
   828 => x"fc80fa51",
   829 => x"96bd2db5",
   830 => x"d408b138",
   831 => x"81ff0bd4",
   832 => x"0cd40853",
   833 => x"81ff0bd4",
   834 => x"0c81ff0b",
   835 => x"d40c81ff",
   836 => x"0bd40c81",
   837 => x"ff0bd40c",
   838 => x"72862a70",
   839 => x"81067656",
   840 => x"51537295",
   841 => x"38b5d408",
   842 => x"549ab904",
   843 => x"73822efe",
   844 => x"e238ff14",
   845 => x"5473feed",
   846 => x"3873b6b8",
   847 => x"0c738b38",
   848 => x"815287fc",
   849 => x"80d05196",
   850 => x"bd2d81ff",
   851 => x"0bd40cd0",
   852 => x"08708f2a",
   853 => x"70810651",
   854 => x"515372f3",
   855 => x"3872d00c",
   856 => x"81ff0bd4",
   857 => x"0c815372",
   858 => x"b5d40c02",
   859 => x"94050d04",
   860 => x"02e8050d",
   861 => x"78558056",
   862 => x"81ff0bd4",
   863 => x"0cd00870",
   864 => x"8f2a7081",
   865 => x"06515153",
   866 => x"72f33882",
   867 => x"810bd00c",
   868 => x"81ff0bd4",
   869 => x"0c775287",
   870 => x"fc80d151",
   871 => x"96bd2d80",
   872 => x"dbc6df54",
   873 => x"b5d40880",
   874 => x"2e8a38b1",
   875 => x"b85185fe",
   876 => x"2d9c8704",
   877 => x"81ff0bd4",
   878 => x"0cd40870",
   879 => x"81ff0651",
   880 => x"537281fe",
   881 => x"2e098106",
   882 => x"9d3880ff",
   883 => x"5395ef2d",
   884 => x"b5d40875",
   885 => x"70840557",
   886 => x"0cff1353",
   887 => x"728025ed",
   888 => x"3881569b",
   889 => x"ec04ff14",
   890 => x"5473c938",
   891 => x"81ff0bd4",
   892 => x"0c81ff0b",
   893 => x"d40cd008",
   894 => x"708f2a70",
   895 => x"81065151",
   896 => x"5372f338",
   897 => x"72d00c75",
   898 => x"b5d40c02",
   899 => x"98050d04",
   900 => x"02e8050d",
   901 => x"77797b58",
   902 => x"55558053",
   903 => x"727625a3",
   904 => x"38747081",
   905 => x"055680f5",
   906 => x"2d747081",
   907 => x"055680f5",
   908 => x"2d525271",
   909 => x"712e8638",
   910 => x"81519cc5",
   911 => x"04811353",
   912 => x"9c9c0480",
   913 => x"5170b5d4",
   914 => x"0c029805",
   915 => x"0d0402ec",
   916 => x"050d7655",
   917 => x"74802ebb",
   918 => x"389a1580",
   919 => x"e02d51a9",
   920 => x"ce2db5d4",
   921 => x"08b5d408",
   922 => x"bcec0cb5",
   923 => x"d4085454",
   924 => x"bcc80880",
   925 => x"2e993894",
   926 => x"1580e02d",
   927 => x"51a9ce2d",
   928 => x"b5d40890",
   929 => x"2b83fff0",
   930 => x"0a067075",
   931 => x"07515372",
   932 => x"bcec0cbc",
   933 => x"ec085372",
   934 => x"802e9938",
   935 => x"bcc008fe",
   936 => x"147129bc",
   937 => x"d40805bc",
   938 => x"f00c7084",
   939 => x"2bbccc0c",
   940 => x"549dda04",
   941 => x"bcd808bc",
   942 => x"ec0cbcdc",
   943 => x"08bcf00c",
   944 => x"bcc80880",
   945 => x"2e8a38bc",
   946 => x"c008842b",
   947 => x"539dd604",
   948 => x"bce00884",
   949 => x"2b5372bc",
   950 => x"cc0c0294",
   951 => x"050d0402",
   952 => x"d8050d80",
   953 => x"0bbcc80c",
   954 => x"845497fd",
   955 => x"2db5d408",
   956 => x"802e9538",
   957 => x"b6bc5280",
   958 => x"519af02d",
   959 => x"b5d40880",
   960 => x"2e8638fe",
   961 => x"549e9004",
   962 => x"ff145473",
   963 => x"8024db38",
   964 => x"738c38b1",
   965 => x"c85185fe",
   966 => x"2d7355a3",
   967 => x"99048056",
   968 => x"810bbcf4",
   969 => x"0c8853b1",
   970 => x"dc52b6f2",
   971 => x"519c902d",
   972 => x"b5d40876",
   973 => x"2e098106",
   974 => x"8738b5d4",
   975 => x"08bcf40c",
   976 => x"8853b1e8",
   977 => x"52b78e51",
   978 => x"9c902db5",
   979 => x"d4088738",
   980 => x"b5d408bc",
   981 => x"f40cbcf4",
   982 => x"08802e80",
   983 => x"f638ba82",
   984 => x"0b80f52d",
   985 => x"ba830b80",
   986 => x"f52d7198",
   987 => x"2b71902b",
   988 => x"07ba840b",
   989 => x"80f52d70",
   990 => x"882b7207",
   991 => x"ba850b80",
   992 => x"f52d7107",
   993 => x"baba0b80",
   994 => x"f52dbabb",
   995 => x"0b80f52d",
   996 => x"71882b07",
   997 => x"535f5452",
   998 => x"5a565755",
   999 => x"7381abaa",
  1000 => x"2e098106",
  1001 => x"8d387551",
  1002 => x"a99e2db5",
  1003 => x"d408569f",
  1004 => x"bf047382",
  1005 => x"d4d52e87",
  1006 => x"38b1f451",
  1007 => x"a08004b6",
  1008 => x"bc527551",
  1009 => x"9af02db5",
  1010 => x"d40855b5",
  1011 => x"d408802e",
  1012 => x"83c73888",
  1013 => x"53b1e852",
  1014 => x"b78e519c",
  1015 => x"902db5d4",
  1016 => x"08893881",
  1017 => x"0bbcc80c",
  1018 => x"a0860488",
  1019 => x"53b1dc52",
  1020 => x"b6f2519c",
  1021 => x"902db5d4",
  1022 => x"08802e8a",
  1023 => x"38b28851",
  1024 => x"85fe2da0",
  1025 => x"e004baba",
  1026 => x"0b80f52d",
  1027 => x"547380d5",
  1028 => x"2e098106",
  1029 => x"80ca38ba",
  1030 => x"bb0b80f5",
  1031 => x"2d547381",
  1032 => x"aa2e0981",
  1033 => x"06ba3880",
  1034 => x"0bb6bc0b",
  1035 => x"80f52d56",
  1036 => x"547481e9",
  1037 => x"2e833881",
  1038 => x"547481eb",
  1039 => x"2e8c3880",
  1040 => x"5573752e",
  1041 => x"09810682",
  1042 => x"d038b6c7",
  1043 => x"0b80f52d",
  1044 => x"55748d38",
  1045 => x"b6c80b80",
  1046 => x"f52d5473",
  1047 => x"822e8638",
  1048 => x"8055a399",
  1049 => x"04b6c90b",
  1050 => x"80f52d70",
  1051 => x"bcc00cff",
  1052 => x"05bcc40c",
  1053 => x"b6ca0b80",
  1054 => x"f52db6cb",
  1055 => x"0b80f52d",
  1056 => x"58760577",
  1057 => x"82802905",
  1058 => x"70bcd00c",
  1059 => x"b6cc0b80",
  1060 => x"f52d70bc",
  1061 => x"e40cbcc8",
  1062 => x"08595758",
  1063 => x"76802e81",
  1064 => x"a3388853",
  1065 => x"b1e852b7",
  1066 => x"8e519c90",
  1067 => x"2db5d408",
  1068 => x"81e738bc",
  1069 => x"c0087084",
  1070 => x"2bbccc0c",
  1071 => x"70bce00c",
  1072 => x"b6e10b80",
  1073 => x"f52db6e0",
  1074 => x"0b80f52d",
  1075 => x"71828029",
  1076 => x"05b6e20b",
  1077 => x"80f52d70",
  1078 => x"84808029",
  1079 => x"12b6e30b",
  1080 => x"80f52d70",
  1081 => x"81800a29",
  1082 => x"1270bce8",
  1083 => x"0cbce408",
  1084 => x"7129bcd0",
  1085 => x"080570bc",
  1086 => x"d40cb6e9",
  1087 => x"0b80f52d",
  1088 => x"b6e80b80",
  1089 => x"f52d7182",
  1090 => x"802905b6",
  1091 => x"ea0b80f5",
  1092 => x"2d708480",
  1093 => x"802912b6",
  1094 => x"eb0b80f5",
  1095 => x"2d70982b",
  1096 => x"81f00a06",
  1097 => x"720570bc",
  1098 => x"d80cfe11",
  1099 => x"7e297705",
  1100 => x"bcdc0c52",
  1101 => x"59524354",
  1102 => x"5e515259",
  1103 => x"525d5759",
  1104 => x"57a39204",
  1105 => x"b6ce0b80",
  1106 => x"f52db6cd",
  1107 => x"0b80f52d",
  1108 => x"71828029",
  1109 => x"0570bccc",
  1110 => x"0c70a029",
  1111 => x"83ff0570",
  1112 => x"892a70bc",
  1113 => x"e00cb6d3",
  1114 => x"0b80f52d",
  1115 => x"b6d20b80",
  1116 => x"f52d7182",
  1117 => x"80290570",
  1118 => x"bce80c7b",
  1119 => x"71291e70",
  1120 => x"bcdc0c7d",
  1121 => x"bcd80c73",
  1122 => x"05bcd40c",
  1123 => x"555e5151",
  1124 => x"55558051",
  1125 => x"9cce2d81",
  1126 => x"5574b5d4",
  1127 => x"0c02a805",
  1128 => x"0d0402ec",
  1129 => x"050d7670",
  1130 => x"872c7180",
  1131 => x"ff065556",
  1132 => x"54bcc808",
  1133 => x"8a387388",
  1134 => x"2c7481ff",
  1135 => x"065455b6",
  1136 => x"bc52bcd0",
  1137 => x"0815519a",
  1138 => x"f02db5d4",
  1139 => x"0854b5d4",
  1140 => x"08802eb3",
  1141 => x"38bcc808",
  1142 => x"802e9838",
  1143 => x"728429b6",
  1144 => x"bc057008",
  1145 => x"5253a99e",
  1146 => x"2db5d408",
  1147 => x"f00a0653",
  1148 => x"a4850472",
  1149 => x"10b6bc05",
  1150 => x"7080e02d",
  1151 => x"5253a9ce",
  1152 => x"2db5d408",
  1153 => x"53725473",
  1154 => x"b5d40c02",
  1155 => x"94050d04",
  1156 => x"02e0050d",
  1157 => x"7970842c",
  1158 => x"bcf00805",
  1159 => x"718f0652",
  1160 => x"55537289",
  1161 => x"38b6bc52",
  1162 => x"73519af0",
  1163 => x"2d72a029",
  1164 => x"b6bc0554",
  1165 => x"807480f5",
  1166 => x"2d565374",
  1167 => x"732e8338",
  1168 => x"81537481",
  1169 => x"e52e81ef",
  1170 => x"38817074",
  1171 => x"06545872",
  1172 => x"802e81e3",
  1173 => x"388b1480",
  1174 => x"f52d7083",
  1175 => x"2a790658",
  1176 => x"56769838",
  1177 => x"b4980853",
  1178 => x"72883872",
  1179 => x"babc0b81",
  1180 => x"b72d76b4",
  1181 => x"980c7353",
  1182 => x"a6b90475",
  1183 => x"8f2e0981",
  1184 => x"0681b438",
  1185 => x"749f068d",
  1186 => x"29baaf11",
  1187 => x"51538114",
  1188 => x"80f52d73",
  1189 => x"70810555",
  1190 => x"81b72d83",
  1191 => x"1480f52d",
  1192 => x"73708105",
  1193 => x"5581b72d",
  1194 => x"851480f5",
  1195 => x"2d737081",
  1196 => x"055581b7",
  1197 => x"2d871480",
  1198 => x"f52d7370",
  1199 => x"81055581",
  1200 => x"b72d8914",
  1201 => x"80f52d73",
  1202 => x"70810555",
  1203 => x"81b72d8e",
  1204 => x"1480f52d",
  1205 => x"73708105",
  1206 => x"5581b72d",
  1207 => x"901480f5",
  1208 => x"2d737081",
  1209 => x"055581b7",
  1210 => x"2d921480",
  1211 => x"f52d7370",
  1212 => x"81055581",
  1213 => x"b72d9414",
  1214 => x"80f52d73",
  1215 => x"70810555",
  1216 => x"81b72d96",
  1217 => x"1480f52d",
  1218 => x"73708105",
  1219 => x"5581b72d",
  1220 => x"981480f5",
  1221 => x"2d737081",
  1222 => x"055581b7",
  1223 => x"2d9c1480",
  1224 => x"f52d7370",
  1225 => x"81055581",
  1226 => x"b72d9e14",
  1227 => x"80f52d73",
  1228 => x"81b72d77",
  1229 => x"b4980c80",
  1230 => x"5372b5d4",
  1231 => x"0c02a005",
  1232 => x"0d0402cc",
  1233 => x"050d7e60",
  1234 => x"5e5a800b",
  1235 => x"bcec08bc",
  1236 => x"f008595c",
  1237 => x"568058bc",
  1238 => x"cc08782e",
  1239 => x"81ae3877",
  1240 => x"8f06a017",
  1241 => x"5754738f",
  1242 => x"38b6bc52",
  1243 => x"76518117",
  1244 => x"579af02d",
  1245 => x"b6bc5680",
  1246 => x"7680f52d",
  1247 => x"56547474",
  1248 => x"2e833881",
  1249 => x"547481e5",
  1250 => x"2e80f638",
  1251 => x"81707506",
  1252 => x"555c7380",
  1253 => x"2e80ea38",
  1254 => x"8b1680f5",
  1255 => x"2d980659",
  1256 => x"7880de38",
  1257 => x"8b537c52",
  1258 => x"75519c90",
  1259 => x"2db5d408",
  1260 => x"80cf389c",
  1261 => x"160851a9",
  1262 => x"9e2db5d4",
  1263 => x"08841b0c",
  1264 => x"9a1680e0",
  1265 => x"2d51a9ce",
  1266 => x"2db5d408",
  1267 => x"b5d40888",
  1268 => x"1c0cb5d4",
  1269 => x"085555bc",
  1270 => x"c808802e",
  1271 => x"98389416",
  1272 => x"80e02d51",
  1273 => x"a9ce2db5",
  1274 => x"d408902b",
  1275 => x"83fff00a",
  1276 => x"06701651",
  1277 => x"5473881b",
  1278 => x"0c787a0c",
  1279 => x"7b54a8c2",
  1280 => x"04811858",
  1281 => x"bccc0878",
  1282 => x"26fed438",
  1283 => x"bcc80880",
  1284 => x"2eae387a",
  1285 => x"51a3a22d",
  1286 => x"b5d408b5",
  1287 => x"d40880ff",
  1288 => x"fffff806",
  1289 => x"555b7380",
  1290 => x"fffffff8",
  1291 => x"2e9238b5",
  1292 => x"d408fe05",
  1293 => x"bcc00829",
  1294 => x"bcd40805",
  1295 => x"57a6d504",
  1296 => x"805473b5",
  1297 => x"d40c02b4",
  1298 => x"050d0402",
  1299 => x"f4050d74",
  1300 => x"70088105",
  1301 => x"710c7008",
  1302 => x"bcc40806",
  1303 => x"5353718e",
  1304 => x"38881308",
  1305 => x"51a3a22d",
  1306 => x"b5d40888",
  1307 => x"140c810b",
  1308 => x"b5d40c02",
  1309 => x"8c050d04",
  1310 => x"02f0050d",
  1311 => x"75881108",
  1312 => x"fe05bcc0",
  1313 => x"0829bcd4",
  1314 => x"08117208",
  1315 => x"bcc40806",
  1316 => x"05795553",
  1317 => x"54549af0",
  1318 => x"2d029005",
  1319 => x"0d0402f4",
  1320 => x"050d7470",
  1321 => x"882a83fe",
  1322 => x"80067072",
  1323 => x"982a0772",
  1324 => x"882b87fc",
  1325 => x"80800673",
  1326 => x"982b81f0",
  1327 => x"0a067173",
  1328 => x"0707b5d4",
  1329 => x"0c565153",
  1330 => x"51028c05",
  1331 => x"0d0402f8",
  1332 => x"050d028e",
  1333 => x"0580f52d",
  1334 => x"74882b07",
  1335 => x"7083ffff",
  1336 => x"06b5d40c",
  1337 => x"51028805",
  1338 => x"0d0402f4",
  1339 => x"050d7476",
  1340 => x"78535452",
  1341 => x"80712597",
  1342 => x"38727081",
  1343 => x"055480f5",
  1344 => x"2d727081",
  1345 => x"055481b7",
  1346 => x"2dff1151",
  1347 => x"70eb3880",
  1348 => x"7281b72d",
  1349 => x"028c050d",
  1350 => x"0402e805",
  1351 => x"0d775680",
  1352 => x"70565473",
  1353 => x"7624b138",
  1354 => x"bccc0874",
  1355 => x"2eaa3873",
  1356 => x"51a4902d",
  1357 => x"b5d408b5",
  1358 => x"d4080981",
  1359 => x"0570b5d4",
  1360 => x"08079f2a",
  1361 => x"77058117",
  1362 => x"57575353",
  1363 => x"74762488",
  1364 => x"38bccc08",
  1365 => x"7426d838",
  1366 => x"72b5d40c",
  1367 => x"0298050d",
  1368 => x"0402f005",
  1369 => x"0db5d008",
  1370 => x"1651aa99",
  1371 => x"2db5d408",
  1372 => x"802e9b38",
  1373 => x"8b53b5d4",
  1374 => x"0852babc",
  1375 => x"51a9ea2d",
  1376 => x"bcf80854",
  1377 => x"73802e86",
  1378 => x"38babc51",
  1379 => x"732d0290",
  1380 => x"050d0402",
  1381 => x"dc050d80",
  1382 => x"705a5574",
  1383 => x"b5d00825",
  1384 => x"af38bccc",
  1385 => x"08752ea8",
  1386 => x"387851a4",
  1387 => x"902db5d4",
  1388 => x"08098105",
  1389 => x"70b5d408",
  1390 => x"079f2a76",
  1391 => x"05811b5b",
  1392 => x"565474b5",
  1393 => x"d0082588",
  1394 => x"38bccc08",
  1395 => x"7926da38",
  1396 => x"805578bc",
  1397 => x"cc082781",
  1398 => x"cd387851",
  1399 => x"a4902db5",
  1400 => x"d408802e",
  1401 => x"81a238b5",
  1402 => x"d4088b05",
  1403 => x"80f52d70",
  1404 => x"842a7081",
  1405 => x"06771078",
  1406 => x"842bbabc",
  1407 => x"0b80f52d",
  1408 => x"5c5c5351",
  1409 => x"55567380",
  1410 => x"2e80c638",
  1411 => x"7416822b",
  1412 => x"adc90bb4",
  1413 => x"a4120c54",
  1414 => x"77753110",
  1415 => x"bcfc1155",
  1416 => x"56907470",
  1417 => x"81055681",
  1418 => x"b72da074",
  1419 => x"81b72d76",
  1420 => x"81ff0681",
  1421 => x"16585473",
  1422 => x"802e8938",
  1423 => x"9c53babc",
  1424 => x"52acca04",
  1425 => x"8b53b5d4",
  1426 => x"0852bcfe",
  1427 => x"1651ad80",
  1428 => x"04741682",
  1429 => x"2baae10b",
  1430 => x"b4a4120c",
  1431 => x"547681ff",
  1432 => x"06811658",
  1433 => x"5473802e",
  1434 => x"89389c53",
  1435 => x"babc52ac",
  1436 => x"f8048b53",
  1437 => x"b5d40852",
  1438 => x"77753110",
  1439 => x"bcfc0551",
  1440 => x"7655a9ea",
  1441 => x"2dad9b04",
  1442 => x"74902975",
  1443 => x"317010bc",
  1444 => x"fc055154",
  1445 => x"b5d40874",
  1446 => x"81b72d81",
  1447 => x"1959748b",
  1448 => x"24a238ab",
  1449 => x"d2047490",
  1450 => x"29753170",
  1451 => x"10bcfc05",
  1452 => x"8c773157",
  1453 => x"51548074",
  1454 => x"81b72d9e",
  1455 => x"14ff1656",
  1456 => x"5474f338",
  1457 => x"02a4050d",
  1458 => x"0402fc05",
  1459 => x"0db5d008",
  1460 => x"1351aa99",
  1461 => x"2db5d408",
  1462 => x"802e8838",
  1463 => x"b5d40851",
  1464 => x"9cce2d80",
  1465 => x"0bb5d00c",
  1466 => x"ab932d8e",
  1467 => x"852d0284",
  1468 => x"050d0402",
  1469 => x"fc050d72",
  1470 => x"5170fd2e",
  1471 => x"ad3870fd",
  1472 => x"248a3870",
  1473 => x"fc2e80c4",
  1474 => x"38aed404",
  1475 => x"70fe2eb1",
  1476 => x"3870ff2e",
  1477 => x"098106bc",
  1478 => x"38b5d008",
  1479 => x"5170802e",
  1480 => x"b338ff11",
  1481 => x"b5d00cae",
  1482 => x"d404b5d0",
  1483 => x"08f00570",
  1484 => x"b5d00c51",
  1485 => x"7080259c",
  1486 => x"38800bb5",
  1487 => x"d00caed4",
  1488 => x"04b5d008",
  1489 => x"8105b5d0",
  1490 => x"0caed404",
  1491 => x"b5d00890",
  1492 => x"05b5d00c",
  1493 => x"ab932d8e",
  1494 => x"852d0284",
  1495 => x"050d0402",
  1496 => x"fc050d80",
  1497 => x"0bb5d00c",
  1498 => x"ab932d8d",
  1499 => x"9c2db5d4",
  1500 => x"08b5c00c",
  1501 => x"b49c518f",
  1502 => x"a02d0284",
  1503 => x"050d0471",
  1504 => x"bcf80c04",
  1505 => x"00ffffff",
  1506 => x"ff00ffff",
  1507 => x"ffff00ff",
  1508 => x"ffffff00",
  1509 => x"20202020",
  1510 => x"203d4b79",
  1511 => x"705a583d",
  1512 => x"20202020",
  1513 => x"00000000",
  1514 => x"20202020",
  1515 => x"20202020",
  1516 => x"20202020",
  1517 => x"20202020",
  1518 => x"00000000",
  1519 => x"52657365",
  1520 => x"74000000",
  1521 => x"4e4d4900",
  1522 => x"43617267",
  1523 => x"61722044",
  1524 => x"6973636f",
  1525 => x"2f43696e",
  1526 => x"74612010",
  1527 => x"00000000",
  1528 => x"45786974",
  1529 => x"00000000",
  1530 => x"4159206d",
  1531 => x"69786572",
  1532 => x"20414342",
  1533 => x"00000000",
  1534 => x"4159206d",
  1535 => x"69786572",
  1536 => x"20414243",
  1537 => x"00000000",
  1538 => x"5363616e",
  1539 => x"6c696e65",
  1540 => x"73204e6f",
  1541 => x"6e650000",
  1542 => x"5363616e",
  1543 => x"6c696e65",
  1544 => x"73204352",
  1545 => x"54203235",
  1546 => x"25000000",
  1547 => x"5363616e",
  1548 => x"6c696e65",
  1549 => x"73204352",
  1550 => x"54203530",
  1551 => x"25000000",
  1552 => x"5363616e",
  1553 => x"6c696e65",
  1554 => x"73204352",
  1555 => x"54203735",
  1556 => x"25000000",
  1557 => x"43617267",
  1558 => x"61204661",
  1559 => x"6c6c6964",
  1560 => x"61000000",
  1561 => x"4f4b0000",
  1562 => x"16200000",
  1563 => x"14200000",
  1564 => x"15200000",
  1565 => x"53442069",
  1566 => x"6e69742e",
  1567 => x"2e2e0a00",
  1568 => x"53442063",
  1569 => x"61726420",
  1570 => x"72657365",
  1571 => x"74206661",
  1572 => x"696c6564",
  1573 => x"210a0000",
  1574 => x"53444843",
  1575 => x"20657272",
  1576 => x"6f72210a",
  1577 => x"00000000",
  1578 => x"57726974",
  1579 => x"65206661",
  1580 => x"696c6564",
  1581 => x"0a000000",
  1582 => x"52656164",
  1583 => x"20666169",
  1584 => x"6c65640a",
  1585 => x"00000000",
  1586 => x"43617264",
  1587 => x"20696e69",
  1588 => x"74206661",
  1589 => x"696c6564",
  1590 => x"0a000000",
  1591 => x"46415431",
  1592 => x"36202020",
  1593 => x"00000000",
  1594 => x"46415433",
  1595 => x"32202020",
  1596 => x"00000000",
  1597 => x"4e6f2070",
  1598 => x"61727469",
  1599 => x"74696f6e",
  1600 => x"20736967",
  1601 => x"0a000000",
  1602 => x"42616420",
  1603 => x"70617274",
  1604 => x"0a000000",
  1605 => x"4261636b",
  1606 => x"00000000",
  1607 => x"00000002",
  1608 => x"00000002",
  1609 => x"00001794",
  1610 => x"00000000",
  1611 => x"00000002",
  1612 => x"000017a8",
  1613 => x"00000000",
  1614 => x"00000002",
  1615 => x"000017bc",
  1616 => x"0000034e",
  1617 => x"00000002",
  1618 => x"000017c4",
  1619 => x"00000379",
  1620 => x"00000003",
  1621 => x"00001994",
  1622 => x"00000004",
  1623 => x"00000003",
  1624 => x"0000198c",
  1625 => x"00000002",
  1626 => x"00000002",
  1627 => x"000017c8",
  1628 => x"0000175f",
  1629 => x"00000002",
  1630 => x"000017e0",
  1631 => x"000006a3",
  1632 => x"00000000",
  1633 => x"00000000",
  1634 => x"00000000",
  1635 => x"000017e8",
  1636 => x"000017f8",
  1637 => x"00001808",
  1638 => x"00001818",
  1639 => x"0000182c",
  1640 => x"00001840",
  1641 => x"00000004",
  1642 => x"00001854",
  1643 => x"000019a4",
  1644 => x"00000004",
  1645 => x"00001864",
  1646 => x"00001920",
  1647 => x"00000000",
  1648 => x"00000000",
  1649 => x"00000000",
  1650 => x"00000000",
  1651 => x"00000000",
  1652 => x"00000000",
  1653 => x"00000000",
  1654 => x"00000000",
  1655 => x"00000000",
  1656 => x"00000000",
  1657 => x"00000000",
  1658 => x"00000000",
  1659 => x"00000000",
  1660 => x"00000000",
  1661 => x"00000000",
  1662 => x"00000000",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00000000",
  1666 => x"00000000",
  1667 => x"00000000",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"00000000",
  1671 => x"00000002",
  1672 => x"00001e7c",
  1673 => x"00001561",
  1674 => x"00000002",
  1675 => x"00001e9a",
  1676 => x"00001561",
  1677 => x"00000002",
  1678 => x"00001eb8",
  1679 => x"00001561",
  1680 => x"00000002",
  1681 => x"00001ed6",
  1682 => x"00001561",
  1683 => x"00000002",
  1684 => x"00001ef4",
  1685 => x"00001561",
  1686 => x"00000002",
  1687 => x"00001f12",
  1688 => x"00001561",
  1689 => x"00000002",
  1690 => x"00001f30",
  1691 => x"00001561",
  1692 => x"00000002",
  1693 => x"00001f4e",
  1694 => x"00001561",
  1695 => x"00000002",
  1696 => x"00001f6c",
  1697 => x"00001561",
  1698 => x"00000002",
  1699 => x"00001f8a",
  1700 => x"00001561",
  1701 => x"00000002",
  1702 => x"00001fa8",
  1703 => x"00001561",
  1704 => x"00000002",
  1705 => x"00001fc6",
  1706 => x"00001561",
  1707 => x"00000002",
  1708 => x"00001fe4",
  1709 => x"00001561",
  1710 => x"00000004",
  1711 => x"00001914",
  1712 => x"00000000",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"000016f3",
  1716 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

